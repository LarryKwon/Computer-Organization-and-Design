module MicroCode #(
	parameter IWIDTH = 26, // control_signal 자리수
	parameter NDEPTH = 256, // control_signal의 가짓수
	parameter AWIDTH = 8 // control_signal의 가짓수를 나타낼 수 있는 index 자리수
) (	
    input wire RSTn,
    input wire[4:0] inst,
    input wire[2:0] stage,
    output wire [IWIDTH-1:0] control_signal // 26자리 배출
);
	//Declare the microcode that will store the control signal
    reg [IWIDTH -1:0] MC [NDEPTH-1:0];

	//Define asynchronous read
    reg [AWIDTH-1:0] index;
    always@(*) begin
        index = {inst[4:0],stage[2:0]};    
    end
	assign control_signal = MC[index];

    initial begin
        //표 작성

        //R-type
        //add
        MC[8'b00000000] <= 11010110000000 // add IF
        MC[8'b00000001] <= 00000000000000 // add ID
        MC[8'b00000010] <= 00000000110000 // add EX
        MC[8'b00000100] <= 00100000000000 // add WB

        //sub
        MC[8'b00001000] <= 11010110000000 // sub IF
        MC[8'b00001001] <= 00000000000000 // sub ID
        MC[8'b00001010] <= 00000000110000 // sub EX
        MC[8'b00001100] <= 00100000000000 // sub WB

        //slt
        MC[8'b00010000] <= 11010110000000 // slt IF
        MC[8'b00010001] <= 00000000000000 // slt ID
        MC[8'b00010010] <= 00000000110000 // slt EX
        MC[8'b00010100] <= 00100000000000 // slt WB

        //sltu
        MC[8'b00011000] <= 11010110000000 // sltu IF
        MC[8'b00011001] <= 00000000000000 // sltu ID
        MC[8'b00011010] <= 00000000100000 // sltu EX
        MC[8'b00011100] <= 00100000000000 // sltu WB

        //xor
        MC[8'b00100000] <= 11010110000000 // xor IF 
        MC[8'b00100001] <= 00000000000000 // xor ID
        MC[8'b00100010] <= 00000000110000 // xor EX
        MC[8'b00100100] <= 00100000000000 // xor WB

        // or
        MC[8'b00101000] <= 11010110000000 // or IF
        MC[8'b00101001] <= 00000000000000 // or ID
        MC[8'b00101010] <= 00000000110000 // or EX
        MC[8'b00101100] <= 00100000000000 // or WB

        //and
        MC[8'b00110000] <= 11010110000000 // and IF
        MC[8'b00110001] <= 00000000000000 // and ID
        MC[8'b00110010] <= 00000000110000 // and EX
        MC[8'b00110100] <= 00100000000000 // and WB

        //sll
        MC[8'b00111000] <= 11010110000000 // sll IF
        MC[8'b00111001] <= 00000000000000 // sll ID
        MC[8'b00111010] <= 00000000110000 // sll EX
        MC[8'b00111100] <= 00100000000000 // sll WB

        //srl
        MC[8'b01000000] <= 11010110000000 // srl IF
        MC[8'b01000001] <= 00000000000000 // srl ID
        MC[8'b01000010] <= 00000000110000 // srl EX
        MC[8'b01000100] <= 00100000000000 // srl WB

        //sra
        MC[8'b01001000] <= 11010110000000 // sra IF
        MC[8'b01001001] <= 00000000000000 // sra ID
        MC[8'b01001010] <= 00000000110000 // sra EX
        MC[8'b01001100] <= 00100000000000 // sra WB

        //I-type
        //add
        MC[8'b01010000] <= 11010110000000 // add IF
        MC[8'b01010001] <= 00000001000000 // add ID
        MC[8'b01010010] <= 00000001110000 // add EX
        MC[8'b01010100] <= 00100001000000 // add WB

        //sub
        MC[8'b01011000] <= 11010110000000 // sub IF
        MC[8'b01011001] <= 00000001000000 // sub ID
        MC[8'b01011010] <= 00000001110000 // sub EX
        MC[8'b01011100] <= 00100001000000 // sub WB

        //slt
        MC[8'b01100000] <= 11010110000000 // slt IF
        MC[8'b01100001] <= 00000001000000 // slt ID
        MC[8'b01100010] <= 00000001110000 // slt EX
        MC[8'b01100100] <= 00100001000000 // slt WB

        //sltu
        MC[8'b01101000] <= 11010110000000 // sltu IF
        MC[8'b01101001] <= 00000001000000 // sltu ID
        MC[8'b01101010] <= 00000001100000 // sltu EX
        MC[8'b01101100] <= 00100001000000 // sltu WB

        //xor
        MC[8'b01110000] <= 11010110000000 // xor IF
        MC[8'b01110001] <= 00000001000000 // xor ID
        MC[8'b01110010] <= 00000001110000 // xor EX
        MC[8'b01110100] <= 00100001000000 // xor WB

        //or
        MC[8'b01111000] <= 11010110000000 // or IF
        MC[8'b01111001] <= 00000001000000 // or ID
        MC[8'b01111010] <= 00000001110000 // or EX
        MC[8'b01111100] <= 00100001000000 // or WB

        //and
        MC[8'b10000000] <= 11010110000000 // and IF
        MC[8'b10000001] <= 00000001000000 // and ID
        MC[8'b10000010] <= 00000001110000 // and EX
        MC[8'b10000100] <= 00100001000000 // and WB

        //sll
        MC[8'b10001000] <= 11010110000000 // sll IF
        MC[8'b10001001] <= 00000001000000 // sll ID
        MC[8'b10001010] <= 00000001110000 // sll EX
        MC[8'b10001100] <= 00100001000000 // sll WB

        //srl
        MC[8'b10010000] <= 11010110000000 // srl IF
        MC[8'b10010001] <= 00000001000000 // srl ID
        MC[8'b10010010] <= 00000001110000 // srl EX
        MC[8'b10010100] <= 00100001000000 // srl WB

        //sra
        MC[8'b10011000] <= 11010110000000 // sra IF
        MC[8'b10011001] <= 00000001000000 // sra ID
        MC[8'b10011010] <= 00000001110000 // sra EX
        MC[8'b10011100] <= 00100001000000 // sra WB

        //L-type
        //LW
        MC[8'10100000] <= 11010110000000// LW IF
        MC[8'10100001] <= 00000001000010// LW ID
        MC[8'10100010] <= 000000011?0010// LW EX
        MC[8'10100011] <= 00000001000010// LW MEM
        MC[8'10100100] <= 00100001000010// LW WB

        //S-type
        //SW
        MC[8'b10101000] <= 11010110000000// SW IF
        MC[8'b10101001] <= 00000001000000// SW ID
        MC[8'b10101010] <= 00000001110000// SW EX
        MC[8'b10101011] <= 00000001000001// SW MEM
        
        //JALR
        MC[8'b10110000] <= 01010001001100// JALR IF
        MC[8'b10110001] <= 00000001001100// JALR ID
        MC[8'b10110010] <= 10000001101100// JALR EX
        MC[8'b10110100] <= 00100110001100// JALR WB
        
        //JAL
        MC[8'b10111000] <= 01010101000000// JALR IF
        MC[8'b10111010] <= 10000101101000// JALR EX
        MC[8'b10111100] <= 00100110001100// JALR WB
                
        //B-type
        //BEQ, BNE, BLT, BGE
        MC[8'b11000000] <= 11010110000000// BXX IF
        MC[8'b11000001] <= 000010011?0000// BXX ID
        MC[8'b11000010] <= 00000000001000// BXX EX

        //BLTU,BGEU
        MC[8'b11001000] <= 11010110000000// BXXU IF
        MC[8'b11001001] <= 000010011?0000// BXXU ID
        MC[8'b11001010] <= 00000000001000// BXXU EX

        //LUI
        MC[8'b11010000] <= 11010110000000// LUI IF
        MC[8'b11010100] <= 00100110000110// LUI WB

        //AUIPC
        MC[8'b11011000] <= 11010110000000// AUIPC IF
        MC[8'b10011010] <= 00000101100000// AUIPC EX
        MC[8'b10011100] <= 00100101000000// AUIPC WB
    end

endmodule